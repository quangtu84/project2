module number (
    input logic enable_i,
    input logic [3:0] number_i,
    input logic [3:0] x_ofs_i,
    input logic [3:0] y_ofs_i,
    output logic number_bit_o
);

    logic [15:0] bit_array [16][16];
    int i,j;
    assign number_bit_o = enable_i ? bit_array[number_i][y_ofs_i][~x_ofs_i] : 0;
    initial begin
        bit_array[0][0]  = 16'b0000_0000_0000_0000;
        bit_array[0][1]  = 16'b0000_1111_1111_0000;
        bit_array[0][2]  = 16'b0000_1111_1111_0000;
        bit_array[0][3]  = 16'b0011_1111_1111_1100;
        bit_array[0][4]  = 16'b0011_1100_0011_1100;
        bit_array[0][5]  = 16'b0011_1100_0011_1100;
        bit_array[0][6]  = 16'b0011_1100_0011_1100;
        bit_array[0][7]  = 16'b0011_1100_0011_1100;
        bit_array[0][8]  = 16'b0011_1100_0011_1100;
        bit_array[0][9]  = 16'b0011_1100_0011_1100;
        bit_array[0][10] = 16'b0011_1100_0011_1100;
        bit_array[0][11] = 16'b0011_1100_0011_1100;
        bit_array[0][12] = 16'b0011_1111_1111_1100;
        bit_array[0][13] = 16'b0000_1111_1111_0000;
        bit_array[0][14] = 16'b0000_1111_1111_0000;
        bit_array[0][15] = 16'b0000_0000_0000_0000;

        bit_array[1][0]  = 16'b0000_0000_0000_0000;
        bit_array[1][1]  = 16'b0000_0011_1100_0000;
        bit_array[1][2]  = 16'b0000_0111_1100_0000;
        bit_array[1][3]  = 16'b0000_1111_1100_0000;
        bit_array[1][4]  = 16'b0001_1111_1100_0000;
        bit_array[1][5]  = 16'b0011_1011_1100_0000;
        bit_array[1][6]  = 16'b0000_0011_1100_0000;
        bit_array[1][7]  = 16'b0000_0011_1100_0000;
        bit_array[1][8]  = 16'b0000_0011_1100_0000;
        bit_array[1][9]  = 16'b0000_0011_1100_0000;
        bit_array[1][10] = 16'b0000_0011_1100_0000;
        bit_array[1][11] = 16'b0000_0011_1100_0000;
        bit_array[1][12] = 16'b0000_0011_1100_0000;
        bit_array[1][13] = 16'b0000_0011_1100_0000;
        bit_array[1][14] = 16'b0000_0011_1100_0000;
        bit_array[1][15] = 16'b0000_0000_0000_0000;

        bit_array[2][0]  = 16'b0000_0000_0000_0000;
        bit_array[2][1]  = 16'b0001_1111_1111_1000;
        bit_array[2][2]  = 16'b0011_1111_1111_1100;
        bit_array[2][3]  = 16'b0011_1111_1111_1100;
        bit_array[2][4]  = 16'b0000_0000_0011_1100;
        bit_array[2][5]  = 16'b0000_0000_0011_1100;
        bit_array[2][6]  = 16'b0001_1111_1111_1100;
        bit_array[2][7]  = 16'b0011_1111_1111_1100;
        bit_array[2][8]  = 16'b0011_1111_1111_1100;
        bit_array[2][9]  = 16'b0011_1111_1111_1000;
        bit_array[2][10] = 16'b0011_1100_0000_0000;
        bit_array[2][11] = 16'b0011_1100_0000_0000;
        bit_array[2][12] = 16'b0011_1111_1111_1100;
        bit_array[2][13] = 16'b0011_1111_1111_1100;
        bit_array[2][14] = 16'b0001_1111_1111_1000;
        bit_array[2][15] = 16'b0000_0000_0000_0000;

        bit_array[3][0]  = 16'b0000_0000_0000_0000;
        bit_array[3][1]  = 16'b0001_1111_1111_1000;
        bit_array[3][2]  = 16'b0011_1111_1111_1100;
        bit_array[3][3]  = 16'b0001_1111_1111_1100;
        bit_array[3][4]  = 16'b0000_0000_0011_1100;
        bit_array[3][5]  = 16'b0000_0000_0011_1100;
        bit_array[3][6]  = 16'b0001_1111_1111_1100;
        bit_array[3][7]  = 16'b0011_1111_1111_1100;
        bit_array[3][8]  = 16'b0011_1111_1111_1100;
        bit_array[3][9]  = 16'b0001_1111_1111_1100;
        bit_array[3][10] = 16'b0000_0000_0011_1100;
        bit_array[3][11] = 16'b0000_0000_0011_1100;
        bit_array[3][12] = 16'b0001_1111_1111_1100;
        bit_array[3][13] = 16'b0011_1111_1111_1100;
        bit_array[3][14] = 16'b0001_1111_1111_1000;
        bit_array[3][15] = 16'b0000_0000_0000_0000;

        bit_array[4][0]  = 16'b0000_0000_0000_0000;
        bit_array[4][1]  = 16'b0001_1100_0011_1100;
        bit_array[4][2]  = 16'b0011_1100_0011_1100;
        bit_array[4][3]  = 16'b0011_1100_0011_1100;
        bit_array[4][4]  = 16'b0011_1100_0011_1100;
        bit_array[4][5]  = 16'b0011_1100_0011_1100;
        bit_array[4][6]  = 16'b0011_1111_1111_1100;
        bit_array[4][7]  = 16'b0011_1111_1111_1100;
        bit_array[4][8]  = 16'b0011_1111_1111_1100;
        bit_array[4][9]  = 16'b0001_1111_1111_1100;
        bit_array[4][10] = 16'b0000_0000_0011_1100;
        bit_array[4][11] = 16'b0000_0000_0011_1100;
        bit_array[4][12] = 16'b0000_0000_0011_1100;
        bit_array[4][13] = 16'b0000_0000_0011_1100;
        bit_array[4][14] = 16'b0000_0000_0011_1100;
        bit_array[4][15] = 16'b0000_0000_0000_0000;

        bit_array[5][0]  = 16'b0000_0000_0000_0000;
        bit_array[5][1]  = 16'b0001_1111_1111_1000;
        bit_array[5][2]  = 16'b0011_1111_1111_1100;
        bit_array[5][3]  = 16'b0011_1111_1111_1100;
        bit_array[5][4]  = 16'b0011_1100_0000_0000;
        bit_array[5][5]  = 16'b0011_1100_0000_0000;
        bit_array[5][6]  = 16'b0011_1111_1111_1000;
        bit_array[5][7]  = 16'b0011_1111_1111_1100;
        bit_array[5][8]  = 16'b0011_1111_1111_1100;
        bit_array[5][9]  = 16'b0001_1111_1111_1100;
        bit_array[5][10] = 16'b0000_0000_0011_1100;
        bit_array[5][11] = 16'b0000_0000_0011_1100;
        bit_array[5][12] = 16'b0001_1111_1111_1100;
        bit_array[5][13] = 16'b0011_1111_1111_1100;
        bit_array[5][14] = 16'b0001_1111_1111_1000;
        bit_array[5][15] = 16'b0000_0000_0000_0000;

        bit_array[6][0]  = 16'b0000_0000_0000_0000;
        bit_array[6][1]  = 16'b0001_1111_1111_1000;
        bit_array[6][2]  = 16'b0011_1111_1111_1100;
        bit_array[6][3]  = 16'b0011_1111_1111_1100;
        bit_array[6][4]  = 16'b0011_1100_0000_0000;
        bit_array[6][5]  = 16'b0011_1100_0000_0000;
        bit_array[6][6]  = 16'b0011_1111_1111_1000;
        bit_array[6][7]  = 16'b0011_1111_1111_1100;
        bit_array[6][8]  = 16'b0011_1111_1111_1100;
        bit_array[6][9]  = 16'b0011_1111_1111_1100;
        bit_array[6][10] = 16'b0011_1100_0011_1100;
        bit_array[6][11] = 16'b0011_1100_0011_1100;
        bit_array[6][12] = 16'b0011_1111_1111_1100;
        bit_array[6][13] = 16'b0011_1111_1111_1100;
        bit_array[6][14] = 16'b0001_1111_1111_1000;
        bit_array[6][15] = 16'b0000_0000_0000_0000;

        bit_array[7][0]  = 16'b0000_0000_0000_0000;
        bit_array[7][1]  = 16'b0001_1111_1111_1000;
        bit_array[7][2]  = 16'b0011_1111_1111_1100;
        bit_array[7][3]  = 16'b0001_1111_1111_1100;
        bit_array[7][4]  = 16'b0000_0000_0011_1100;
        bit_array[7][5]  = 16'b0000_0000_0011_1100;
        bit_array[7][6]  = 16'b0000_0000_0011_1100;
        bit_array[7][7]  = 16'b0000_0000_0011_1100;
        bit_array[7][8]  = 16'b0000_0000_0011_1100;
        bit_array[7][9]  = 16'b0000_0000_0011_1100;
        bit_array[7][10] = 16'b0000_0000_0011_1100;
        bit_array[7][11] = 16'b0000_0000_0011_1100;
        bit_array[7][12] = 16'b0000_0000_0011_1100;
        bit_array[7][13] = 16'b0000_0000_0011_1100;
        bit_array[7][14] = 16'b0000_0000_0011_1100;
        bit_array[7][15] = 16'b0000_0000_0000_0000;

        bit_array[8][0]  = 16'b0000_0000_0000_0000;
        bit_array[8][1]  = 16'b0001_1111_1111_1000;
        bit_array[8][2]  = 16'b0011_1111_1111_1100;
        bit_array[8][3]  = 16'b0011_1111_1111_1100;
        bit_array[8][4]  = 16'b0011_1100_0011_1100;
        bit_array[8][5]  = 16'b0011_1100_0011_1100;
        bit_array[8][6]  = 16'b0011_1111_1111_1100;
        bit_array[8][7]  = 16'b0001_1111_1111_1000;
        bit_array[8][8]  = 16'b0001_1111_1111_1000;
        bit_array[8][9]  = 16'b0011_1111_1111_1100;
        bit_array[8][10] = 16'b0011_1100_0011_1100;
        bit_array[8][11] = 16'b0011_1100_0011_1100;
        bit_array[8][12] = 16'b0011_1111_1111_1100;
        bit_array[8][13] = 16'b0011_1111_1111_1100;
        bit_array[8][14] = 16'b0001_1111_1111_1000;
        bit_array[8][15] = 16'b0000_0000_0000_0000;

        bit_array[9][0]  = 16'b0000_0000_0000_0000;
        bit_array[9][1]  = 16'b0001_1111_1111_1000;
        bit_array[9][2]  = 16'b0011_1111_1111_1100;
        bit_array[9][3]  = 16'b0011_1111_1111_1100;
        bit_array[9][4]  = 16'b0011_1100_0011_1100;
        bit_array[9][5]  = 16'b0011_1100_0011_1100;
        bit_array[9][6]  = 16'b0011_1111_1111_1100;
        bit_array[9][7]  = 16'b0011_1111_1111_1100;
        bit_array[9][8]  = 16'b0011_1111_1111_1100;
        bit_array[9][9]  = 16'b0001_1111_1111_1100;
        bit_array[9][10] = 16'b0000_0000_0011_1100;
        bit_array[9][11] = 16'b0000_0000_0011_1100;
        bit_array[9][12] = 16'b0001_1111_1111_1100;
        bit_array[9][13] = 16'b0011_1111_1111_1100;
        bit_array[9][14] = 16'b0001_1111_1111_1000;
        bit_array[9][15] = 16'b0000_0000_0000_0000;

        for(i = 10; i <= 15; i ++)
            for(j = 0; j <= 15; j ++)
                bit_array[i][j] = 16'b0;

    end
endmodule
