module top #(
    parameter COLOR_BITS = 24
) (
    input logic [3:0] player_1_move_i,
    input logic [3:0] player_2_move_i,
    input logic player_1_shoot_i,
    input logic player_2_shoot_i,
    output logic hsync_no,
    output logic vsync_no,
    //for simulation only
    output logic [9:0] hpos_o,
    output logic [9:0] vpos_o,
    output logic display_enable_o,
    /////////////////////////
    output logic [(COLOR_BITS/3)-1 :0] blue_o,
    output logic [(COLOR_BITS/3)-1 :0] green_o,
    output logic [(COLOR_BITS/3)-1 :0] red_o,
	output logic VGA_clk_o,
    input logic clk_i,
    input logic reset_i
);

    game_top #(
        .COLOR_BITS(COLOR_BITS)
    ) top(
        .*
    );

endmodule
